module addsub32(
  input logic [31:0] i_a,
  input logic [31:0] i_b,
  input logic Cin,
  output logic Cout,
  output logic [31:0] o_s
);

logic [31:0] C;

	always_comb begin
	
		C[0] = Cin;
		
		o_s[0]  = i_a[0]  ^ (i_b[0]  ^ Cin) ^ C[0];
		C[1]  = (i_a[0]  & (i_b[0]  ^ Cin)) | (C[0]  & (i_a[0]  ^ (i_b[0]  ^ Cin)));

		o_s[1]  = i_a[1]  ^ (i_b[1]  ^ Cin) ^ C[1];
		C[2]  = (i_a[1]  & (i_b[1]  ^ Cin)) | (C[1]  & (i_a[1]  ^ (i_b[1]  ^ Cin)));

		o_s[2]  = i_a[2]  ^ (i_b[2]  ^ Cin) ^ C[2];
		C[3]  = (i_a[2]  & (i_b[2]  ^ Cin)) | (C[2]  & (i_a[2]  ^ (i_b[2]  ^ Cin)));

		o_s[3]  = i_a[3]  ^ (i_b[3]  ^ Cin) ^ C[3];
		C[4]  = (i_a[3]  & (i_b[3]  ^ Cin)) | (C[3]  & (i_a[3]  ^ (i_b[3]  ^ Cin)));

		o_s[4]  = i_a[4]  ^ (i_b[4]  ^ Cin) ^ C[4];
		C[5]  = (i_a[4]  & (i_b[4]  ^ Cin)) | (C[4]  & (i_a[4]  ^ (i_b[4]  ^ Cin)));

		o_s[5]  = i_a[5]  ^ (i_b[5]  ^ Cin) ^ C[5];
		C[6]  = (i_a[5]  & (i_b[5]  ^ Cin)) | (C[5]  & (i_a[5]  ^ (i_b[5]  ^ Cin)));

		o_s[6]  = i_a[6]  ^ (i_b[6]  ^ Cin) ^ C[6];
		C[7]  = (i_a[6]  & (i_b[6]  ^ Cin)) | (C[6]  & (i_a[6]  ^ (i_b[6]  ^ Cin)));

		o_s[7]  = i_a[7]  ^ (i_b[7]  ^ Cin) ^ C[7];
		C[8]  = (i_a[7]  & (i_b[7]  ^ Cin)) | (C[7]  & (i_a[7]  ^ (i_b[7]  ^ Cin)));

		o_s[8]  = i_a[8]  ^ (i_b[8]  ^ Cin) ^ C[8];
		C[9]  = (i_a[8]  & (i_b[8]  ^ Cin)) | (C[8]  & (i_a[8]  ^ (i_b[8]  ^ Cin)));

		o_s[9]  = i_a[9]  ^ (i_b[9]  ^ Cin) ^ C[9];
		C[10] = (i_a[9]  & (i_b[9]  ^ Cin)) | (C[9]  & (i_a[9]  ^ (i_b[9]  ^ Cin)));

		o_s[10] = i_a[10] ^ (i_b[10] ^ Cin) ^ C[10];
		C[11] = (i_a[10] & (i_b[10] ^ Cin)) | (C[10] & (i_a[10] ^ (i_b[10] ^ Cin)));

		o_s[11] = i_a[11] ^ (i_b[11] ^ Cin) ^ C[11];
		C[12] = (i_a[11] & (i_b[11] ^ Cin)) | (C[11] & (i_a[11] ^ (i_b[11] ^ Cin)));

		o_s[12] = i_a[12] ^ (i_b[12] ^ Cin) ^ C[12];
		C[13] = (i_a[12] & (i_b[12] ^ Cin)) | (C[12] & (i_a[12] ^ (i_b[12] ^ Cin)));

		o_s[13] = i_a[13] ^ (i_b[13] ^ Cin) ^ C[13];
		C[14] = (i_a[13] & (i_b[13] ^ Cin)) | (C[13] & (i_a[13] ^ (i_b[13] ^ Cin)));

		o_s[14] = i_a[14] ^ (i_b[14] ^ Cin) ^ C[14];
		C[15] = (i_a[14] & (i_b[14] ^ Cin)) | (C[14] & (i_a[14] ^ (i_b[14] ^ Cin)));

		o_s[15] = i_a[15] ^ (i_b[15] ^ Cin) ^ C[15];
		C[16] = (i_a[15] & (i_b[15] ^ Cin)) | (C[15] & (i_a[15] ^ (i_b[15] ^ Cin)));

		o_s[16] = i_a[16] ^ (i_b[16] ^ Cin) ^ C[16];
		C[17] = (i_a[16] & (i_b[16] ^ Cin)) | (C[16] & (i_a[16] ^ (i_b[16] ^ Cin)));

		o_s[17] = i_a[17] ^ (i_b[17] ^ Cin) ^ C[17];
		C[18] = (i_a[17] & (i_b[17] ^ Cin)) | (C[17] & (i_a[17] ^ (i_b[17] ^ Cin)));

		o_s[18] = i_a[18] ^ (i_b[18] ^ Cin) ^ C[18];
		C[19] = (i_a[18] & (i_b[18] ^ Cin)) | (C[18] & (i_a[18] ^ (i_b[18] ^ Cin)));

		o_s[19] = i_a[19] ^ (i_b[19] ^ Cin) ^ C[19];
		C[20] = (i_a[19] & (i_b[19] ^ Cin)) | (C[19] & (i_a[19] ^ (i_b[19] ^ Cin)));

		o_s[20] = i_a[20] ^ (i_b[20] ^ Cin) ^ C[20];
		C[21] = (i_a[20] & (i_b[20] ^ Cin)) | (C[20] & (i_a[20] ^ (i_b[20] ^ Cin)));

		o_s[21] = i_a[21] ^ (i_b[21] ^ Cin) ^ C[21];
		C[22] = (i_a[21] & (i_b[21] ^ Cin)) | (C[21] & (i_a[21] ^ (i_b[21] ^ Cin)));

		o_s[22] = i_a[22] ^ (i_b[22] ^ Cin) ^ C[22];
		C[23] = (i_a[22] & (i_b[22] ^ Cin)) | (C[22] & (i_a[22] ^ (i_b[22] ^ Cin)));

		o_s[23] = i_a[23] ^ (i_b[23] ^ Cin) ^ C[23];
		C[24] = (i_a[23] & (i_b[23] ^ Cin)) | (C[23] & (i_a[23] ^ (i_b[23] ^ Cin)));

		o_s[24] = i_a[24] ^ (i_b[24] ^ Cin) ^ C[24];
		C[25] = (i_a[24] & (i_b[24] ^ Cin)) | (C[24] & (i_a[24] ^ (i_b[24] ^ Cin)));

		o_s[25] = i_a[25] ^ (i_b[25] ^ Cin) ^ C[25];
		C[26] = (i_a[25] & (i_b[25] ^ Cin)) | (C[25] & (i_a[25] ^ (i_b[25] ^ Cin)));

		o_s[26] = i_a[26] ^ (i_b[26] ^ Cin) ^ C[26];
		C[27] = (i_a[26] & (i_b[26] ^ Cin)) | (C[26] & (i_a[26] ^ (i_b[26] ^ Cin)));

		o_s[27] = i_a[27] ^ (i_b[27] ^ Cin) ^ C[27];
		C[28] = (i_a[27] & (i_b[27] ^ Cin)) | (C[27] & (i_a[27] ^ (i_b[27] ^ Cin)));

		o_s[28] = i_a[28] ^ (i_b[28] ^ Cin) ^ C[28];
		C[29] = (i_a[28] & (i_b[28] ^ Cin)) | (C[28] & (i_a[28] ^ (i_b[28] ^ Cin)));

		o_s[29] = i_a[29] ^ (i_b[29] ^ Cin) ^ C[29];
		C[30] = (i_a[29] & (i_b[29] ^ Cin)) | (C[29] & (i_a[29] ^ (i_b[29] ^ Cin)));

		o_s[30] = i_a[30] ^ (i_b[30] ^ Cin) ^ C[30];
		C[31] = (i_a[30] & (i_b[30] ^ Cin)) | (C[30] & (i_a[30] ^ (i_b[30] ^ Cin)));

		o_s[31] = i_a[31] ^ (i_b[31] ^ Cin) ^ C[31];
		Cout = (i_a[31] & (i_b[31] ^ Cin)) | (C[31] & (i_a[31] ^ (i_b[31] ^ Cin)));

	end
	
endmodule